library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity tb_mainCircuit is
--  Port ( );
end tb_mainCircuit;

architecture Behavioral of tb_mainCircuit is

begin


end Behavioral;
